#bin/sh
sftp -p 10021 plaza01@plaza.ekankyo21.com
#pass: P56a-MN4df
#https://plaza.ekankyo21.com/
#ID： plaza
#Pass： Pass26za